module resErr(
        
    );
endmodule
